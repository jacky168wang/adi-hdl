
/*
//
//  Module:       cp_removal
//
//  Description:  cyclic prefix removal to FFT size.
//
//  Maintainer:   Royce Ai Yu Pan
//
//  Revision:     0.30
//
//  Change Log:   0.10 2018/01/30, initial draft.
//                0.20 2018/02/23, symbol data always enable supported.
//                0.30 2018/05/26, zip-zap trigger supported.
//                0.40 2018/12/10, blocfifo_inst added.
//
*/

`timescale 1ns/100ps

module cp_removal #(
  
  parameter FFT_SIZE = 4096,                    // FFT size
  parameter CP_LEN1 = 352,                      // long cp length
  parameter CP_LEN2 = 288,                      // short cp length
  parameter BLOCK_QTY = 2,                      // block quantity
  parameter BLOC_ADDR_WIDTH = 2,                // block address bit width, able to represent maximum BLOCK_QTY required.  
  parameter OFFS_ADDR_WIDTH = 13,               // offset address bit width
  parameter WORD_ADDR_WIDTH = 14,               // word address bit width  
  parameter INDX_WIDTH_RD = 13,                 // output data index bit width
  parameter DIN_READY_ADV = 1'b1,               // input ready assert advance
  parameter BLOC_FULL_THRES = 0,                // block full threshold
  parameter BLOC_EMPTY_THRES = 0,               // block empty threshold
  parameter READ_DURING_WRITE = 1'b1,           // read during write
  parameter DOUT_READY_REQ = 1                  // output ready as request  
        
  ) (
  
  input clk_wr,                                 // write clock, posedge active
  input clk_rd,                                 // read clock, posedge active
  input rst_n,                                  // reset, low active
    
  input din_restart,                            // input data restart                                                                                                                                                                                                                                                                                                                                                                                                                                                          
  input din_valid,                              // input data valid
  input din_sop,                                // input data sop
  input din_eop,                                // input data eop  
  input [15:0] din_real,                        // input data real
  input [15:0] din_imag,                        // input data imaginary
  input [1:0] dout_enable,                      // output enable, bit 0 for dout_real and bit 1 for dout_imag.
  input dmem_always,                            // symbol data always enable. not latched, shall not change while operating.
  input [1:0] din_ante,                         // input din_ante  
  input [3:0] din_symbol,                       // input symbol index
  input [7:0] din_slot,                         // input slot index  
  input [9:0] din_frame,                        // input frame index 
  input long_cp,                                // long cyclic prefix
  input dout_trigger,                           // output trigger
  input dout_sync,                              // output sync with long cyclic prefix
  input dout_drop,                              // output data drop
  input dout_repeat,                            // output data repeat
  input dout_ready,                             // output ready        
 
  output din_ready,                             // input ready
  output sop_wr_m,                              // memory write start of packet
  output eop_wr_m,                              // memory write end of packet
  output dmem_valid,                            // symbol data valid
  output dout_sop,                              // output start of packet
  output dout_eop,                              // output end of packet
  output dout_valid,                            // output data valid
  output [15:0] dout_real,                      // output data real
  output [15:0] dout_imag,                      // output data imaginary 
  output [1:0]  dout_ante,                      // dout_ante index
  output [1:0]  dout_ante_pre,                  // predictive dout_ante
  output [3:0]  dout_symbol,                    // output symbol index
  output [3:0]  dout_symbol_pre,                // predictive output symbol index
  output [7:0]  dout_slot,                      // output slot index
  output [7:0]  dout_slot_pre,                  // predictive output slot index
  output [9:0]  dout_frame,                     // output frame index
  output [9:0]  dout_frame_pre,                 // predictive output frame index                
  output [INDX_WIDTH_RD-1:0] dout_index,        // output data index
  output [INDX_WIDTH_RD-1:0] din_index,         // input data index
  output reg [31:0] overflow_cnt,               // block overflow count
  output [WORD_ADDR_WIDTH:0] word_used_drw,     // word used quantity during write, minimum 0 and maximum 'BLOCK_LEN_WR * BLOCK_QTY'.
  output [BLOC_ADDR_WIDTH-1:0] bloc_used,       // block used quantity, minimum 0 and maximum BLOCK_QTY.
  output bloc_full,                             // block full
  output bloc_empty                             // block empty  
              
  );
  
  localparam LATENCY_RD = 2;  
  
  wire dmem_restart;
  wire din_sop_r;
  wire din_eop_r;
  wire eop_rd_m;
  wire en_wr_m;    
  wire [BLOC_ADDR_WIDTH-1:0] bloc_used_rd;
  wire [BLOC_ADDR_WIDTH-1:0] bloc_addr_wr_m;
  wire [BLOC_ADDR_WIDTH-1:0] bloc_addr_rd_m; 
  reg  [BLOC_ADDR_WIDTH-1:0] bloc_addr_rd_m_r0; 
  reg  [BLOC_ADDR_WIDTH-1:0] bloc_addr_rd_m_r1;   
  wire [BLOC_ADDR_WIDTH-1:0] bloc_addr_rd_m_pre;
  wire [WORD_ADDR_WIDTH-1:0] word_addr_wr_m;
  wire [WORD_ADDR_WIDTH-2:0] word_addr_rd_m;  
  wire [15:0] data_real;   
  wire [15:0] data_imag;   
  wire [15:0] data_real_wr_m;
  wire [15:0] data_imag_wr_m;
  wire [15:0] dmem_real;
  wire [15:0] dmem_imag; 
  reg  [15:0] dmem_real_r;
  reg  [15:0] dmem_imag_r;    
  wire dmem_drop;
  wire dmem_request;  
  reg  [1:0]dmem_enable;
  reg  dout_request;
  wire dmem_sop;
  wire dmem_eop;
  wire dout_sop_s;      
  wire dout_valid_s;    
  reg  [INDX_WIDTH_RD-1:0] dmem_index;
  reg  [INDX_WIDTH_RD-1:0] dmem_index_cc[2:1];   
  reg  bloc_full_r;    
  wire [1:0] symbol_sop;
  wire [1:0] symbol_eop;
  wire trigger_start;
  reg  dout_trigger_dly;
  reg  zip_zap;  
  reg  [1:0] symbol_long_cp;
  reg  [1:0] symbol_valid;
  reg  [INDX_WIDTH_RD-1:0] symbol_index [1:0];
  reg  [1:0] ante_list   [BLOCK_QTY-1:0];   
  reg  [3:0] symbol_list [BLOCK_QTY-1:0];
  reg  [7:0] slot_list   [BLOCK_QTY-1:0];
  reg  [9:0] frame_list  [BLOCK_QTY-1:0]; 
  
  assign bloc_full = bloc_used == BLOCK_QTY;   
  assign dmem_drop = 1'b0;
  assign dmem_restart = bloc_full | bloc_full_r;  
  assign dmem_request = DOUT_READY_REQ ? dout_ready : dout_request;           
  assign dmem_valid = dmem_enable[0] & symbol_index[0] >= (symbol_long_cp[0] ? CP_LEN1 : CP_LEN2) & symbol_index[0] <= (symbol_long_cp[0] ? CP_LEN1 : CP_LEN2) + FFT_SIZE - 1
                    | dmem_enable[1] & symbol_index[1] >= (symbol_long_cp[1] ? CP_LEN1 : CP_LEN2) & symbol_index[1] <= (symbol_long_cp[1] ? CP_LEN1 : CP_LEN2) + FFT_SIZE - 1;
  assign data_real = (dmem_valid | dmem_always & |symbol_valid) & dout_enable[0] ? din_real : 16'd0;
  assign data_imag = (dmem_valid | dmem_always & |symbol_valid) & dout_enable[1] ? din_imag : 16'd0;
  assign dmem_sop = dmem_valid & (symbol_sop[0] | symbol_sop[1]);
  assign dmem_eop = dmem_valid & (symbol_eop[0] | symbol_eop[1]);
  assign symbol_sop[0] = symbol_index[0] == (symbol_long_cp[0] ? CP_LEN1 : CP_LEN2);
  assign symbol_sop[1] = symbol_index[1] == (symbol_long_cp[1] ? CP_LEN1 : CP_LEN2);
  assign symbol_eop[0] = symbol_index[0] == (symbol_long_cp[0] ? CP_LEN1 : CP_LEN2) + FFT_SIZE - 1;
  assign symbol_eop[1] = symbol_index[1] == (symbol_long_cp[1] ? CP_LEN1 : CP_LEN2) + FFT_SIZE - 1;
  assign trigger_start = dout_trigger & ~dout_trigger_dly;
  assign din_ready = DIN_READY_ADV ? trigger_start | symbol_valid[0] & ~symbol_eop[0] | symbol_valid[1] & ~symbol_eop[1] : |symbol_valid;
  assign din_sop_r = symbol_valid[0] & symbol_index[0] == 0 | symbol_valid[1] & symbol_index[1] == 0;
  assign din_eop_r = symbol_eop[0] | symbol_eop[1];
  assign din_index = zip_zap ? symbol_index[1] : symbol_index[0];   
  assign dout_sop = dout_sop_s;
  assign dout_valid = dout_valid_s;             
  assign dout_real = dout_valid_s & dout_enable[0] ? dmem_real_r : 15'd0;      
  assign dout_imag = dout_valid_s & dout_enable[1] ? dmem_imag_r: 15'd0; 
  assign bloc_addr_rd_m_pre = bloc_addr_rd_m_r1 == BLOCK_QTY - 1 ? 0 : bloc_addr_rd_m_r1 + 1'b1;         
  assign dout_ante = ante_list[bloc_addr_rd_m_r1];   
  assign dout_symbol = symbol_list[bloc_addr_rd_m_r1];
  assign dout_slot = slot_list[bloc_addr_rd_m_r1];
  assign dout_frame = frame_list[bloc_addr_rd_m_r1];
  assign dout_ante_pre = ante_list[bloc_addr_rd_m_pre];    
  assign dout_symbol_pre = symbol_list[bloc_addr_rd_m_pre];
  assign dout_slot_pre = slot_list[bloc_addr_rd_m_pre];
  assign dout_frame_pre = frame_list[bloc_addr_rd_m_pre];  
  
  integer i;
  
  always @(posedge clk_wr or negedge rst_n) begin
    for(i = 0; i < BLOCK_QTY; i = i + 1) begin
      if(! rst_n) begin
      	ante_list[i]   <= 2'd0;      	        
        symbol_list[i] <= 4'd0;
        slot_list[i]   <= 8'd0;
        frame_list[i]  <= 10'd0;
      end
      else if(sop_wr_m & bloc_addr_wr_m == i) begin
      	ante_list[i]   <= din_ante;      	       
        symbol_list[i] <= din_symbol;
        slot_list[i]   <= din_slot;
        frame_list[i]  <= din_frame;
      end
    end
  end  
  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      bloc_full_r <= 1'b1;
    end
    else if(bloc_full) begin
      bloc_full_r <= 1'b1;
    end
    else if(din_sop_r & din_valid) begin
      bloc_full_r <= 1'b0;
    end
  end
  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      overflow_cnt <= 32'd0;
    end
    else if(dmem_eop & dmem_valid & dmem_restart) begin
      overflow_cnt <= overflow_cnt + 1'b1;
    end
  end  

  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      dmem_index <= 0;
    end
    else if(dmem_valid) begin
      dmem_index <= dmem_eop ? 0 : dmem_index + 1'b1;
    end
  end
  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      zip_zap <= 1'b0;
    end
    else if(trigger_start) begin
      zip_zap <= ~zip_zap;
    end
  end
  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      symbol_long_cp[0] <= 1'b0;
    end
    else if(trigger_start & zip_zap) begin
      symbol_long_cp[0] <= long_cp;
    end
  end
  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      symbol_long_cp[1] <= 1'b0;
    end
    else if(trigger_start & ~zip_zap) begin
      symbol_long_cp[1] <= long_cp;
    end
  end
  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      symbol_valid[0] <= 1'b0;
    end
    else if(trigger_start & zip_zap) begin
      symbol_valid[0] <= 1'b1;
    end
    else if(symbol_eop[0]) begin
      symbol_valid[0] <= 1'b0;
    end
  end
  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      symbol_valid[1] <= 1'b0;
    end
    else if(trigger_start & ~zip_zap) begin
      symbol_valid[1] <= 1'b1;
    end
    else if(symbol_eop[1]) begin
      symbol_valid[1] <= 1'b0;
    end
  end
  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      symbol_index[0] <= 0;
    end
    else if(trigger_start & zip_zap | symbol_eop[0]) begin
      symbol_index[0] <= 0;
    end
    else if(symbol_valid[0]) begin
      symbol_index[0] <= symbol_index[0] + 1'b1;
    end
  end
  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      symbol_index[1] <= 0;
    end
    else if(trigger_start & ~zip_zap | symbol_eop[1]) begin
      symbol_index[1] <= 0;
    end
    else if(symbol_valid[1]) begin
      symbol_index[1] <= symbol_index[1] + 1'b1;
    end
  end
  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      dmem_enable[0] <= 1'b0;
    end
    else if(trigger_start & zip_zap & dmem_enable[1]) begin
      dmem_enable[0] <= din_valid & ~bloc_full;
    end
    else if(trigger_start & zip_zap & (long_cp | ~dout_sync)) begin
      dmem_enable[0] <= din_valid & ~bloc_full;
    end
    else if(symbol_eop[0]) begin
      dmem_enable[0] <= 1'b0;
    end
  end
  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      dmem_enable[1] <= 1'b0;
    end
    else if(trigger_start & ~zip_zap & dmem_enable[0]) begin
      dmem_enable[1] <= din_valid & ~bloc_full;
    end
    else if(trigger_start & ~zip_zap & (long_cp | ~dout_sync)) begin
      dmem_enable[1] <= din_valid & ~bloc_full;
    end
    else if(symbol_eop[1]) begin
      dmem_enable[1] <= 1'b0;
    end
  end
  
  always @(posedge clk_rd or negedge rst_n) begin             
    if(! rst_n) begin                                         
      dmem_index_cc[1] <= 0;  
      dmem_index_cc[2] <= 0;                                            
    end  
    else begin
    	dmem_index_cc[1] <= dmem_index ;    
    	dmem_index_cc[2] <= dmem_index_cc[1];  
    end
  end   
  
  always @(posedge clk_rd or negedge rst_n) begin
    if(! rst_n) begin
      dout_request <= 1'b0;
    end           
    else if(~dout_request & ~dout_valid_s | eop_rd_m) begin
      dout_request <= ( (bloc_used_rd == 0 & dmem_index_cc[2] >= FFT_SIZE/2 + 1) | bloc_used_rd>=1 ) & dout_ready ;
    end
  end 
  
//  always @(posedge clk_rd or negedge rst_n) begin
//   if(! rst_n) begin
//     dout_request <= 1'b0;
//   end
//   else if(eop_rd_m) begin
//     dout_request <= (bloc_used_rd >= 2 | bloc_used_rd >= 1 & dout_repeat) & dout_ready ;
//   end
//   else if(~dout_request & ~dout_valid_s) begin
//     dout_request <= bloc_used_rd >= 1 & dout_ready ;
//   end
// end 

  
  always @(posedge clk_wr or negedge rst_n) begin
    if(! rst_n) begin
      dout_trigger_dly <= 1'b1;
    end
    else begin
      dout_trigger_dly <= dout_trigger;
    end
  end
  
  always @(posedge clk_rd or negedge rst_n) begin                        
    if(! rst_n) begin                                                    
      dmem_real_r <= 0;
      dmem_imag_r <= 0;                                           
    end                                                                  
    else begin                                                           
      dmem_real_r <= dmem_real;     
      dmem_imag_r <= dmem_imag;   
    end                                                                  
  end  
  
  always @(posedge clk_rd or negedge rst_n) begin                     
    if(! rst_n) begin                                                 
      bloc_addr_rd_m_r0 <= 0;                                               
      bloc_addr_rd_m_r1 <= 0;                                               
    end                                                               
    else begin                                                        
      bloc_addr_rd_m_r0 <= bloc_addr_rd_m;                                       
      bloc_addr_rd_m_r1 <= bloc_addr_rd_m_r0;                                       
    end                                                               
  end                                                                 
  
  util_blocfifo #(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
    .DATA_WIDTH_WR(32),                           // write data bit width                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  
    .DATA_WIDTH_RD(32),                           // read data bit width                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
    .BLOCK_LEN_WR(FFT_SIZE),                      // write data block length                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               
    .BLOCK_LEN_RD(FFT_SIZE),                      // read data block length                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                
    .BLOCK_QTY(BLOCK_QTY),                        // block quantity                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        
    .BLOC_ADDR_WIDTH(BLOC_ADDR_WIDTH),            // block address bit width, able to represent maximum BLOCK_QTY required.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                
    .OFFS_ADDR_WIDTH(OFFS_ADDR_WIDTH),            // offset address bit width, able to represent maximum 'BLOCK_LEN_WR - 1' and 'BLOCK_LEN_RD - 1' required.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               
    .WORD_ADDR_WIDTH(WORD_ADDR_WIDTH),            // word address bit width                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                
    .INDX_WIDTH_RD(INDX_WIDTH_RD),                // output data index bit width                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           
    .SEGMENT_QTY(1),                              // read data segment quantity, minimum 1 required.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       
    .SEGM_ADDR_WIDTH(1),                          // segment address bit width, able to represent maximum 'SEGMENT_QTY - 1' required.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      
    .PROFILE_QTY(1),                              // segment profile quantity, minimum 1 required.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
    .PROF_SEL_WIDTH(1),                           // segment profile select bit width, able to represent maximum 'PROFILE_QTY - 1' required.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               
    .SEGM_START('{'{0}}),                         // segment start offset address                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           
    .SEGM_END('{'{FFT_SIZE-1}}),                  // segment end offset address                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  
    .SEGM_STEP('{'{1}}),                          // segment offset address step                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       
    .BLOC_FULL_THRES(BLOC_FULL_THRES),            // block full threshold                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  
    .BLOC_EMPTY_THRES(BLOC_EMPTY_THRES),          // block empty threshold                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 
    .READ_DURING_WRITE(READ_DURING_WRITE),        // read during write                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
    .LATENCY_RD(LATENCY_RD)                       // read data latency, minimum 1.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
  ) blocfifo_inst (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        
    .clk_wr(clk_wr),                              // write clock, posedge active                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           
    .clk_rd(clk_rd),                              // read clock, posedge active                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            
    .rst_n(rst_n),                                // reset, low active                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     
    .mode_sel(dout_repeat),                       // block mode select, '0' - block clear, '1' - block hold.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               
    .din_restart(dmem_restart | din_restart),     // input data restart                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    
    .din_valid(dmem_valid),                       // input data valid                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      
    .din_data({data_imag, data_real}),            // input data                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            
    .prof_sel(1'b0),                              // segment profile select, '0' - profile 0, '1' - profile 1, ...                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
    .dout_drop(dmem_drop | dout_drop),            // output data drop                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      
    .dout_restart(1'b0),                          // output data restart                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
    .dout_request(dmem_request),                  // output data request                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                
    .din_ready(),                                 // input ready                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
    .dout_sop(dout_sop_s),                        // output start of packet                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
    .dout_eop(dout_eop),                          // output end of packet                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                
    .dout_valid(dout_valid_s),                    // output data valid                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
    .dout_data(),                                 // output data                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
    .dout_index(dout_index),                      // output data index                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
    .word_used_drw_wr(),                          // word used quantity during write, on write clock, minimum 0 and maximum 'BLOCK_LEN_WR * BLOCK_QTY'.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  
    .word_used_drw_rd(word_used_drw),             // word used quantity during write, on read clock, minimum 0 and maximum 'BLOCK_LEN_WR * BLOCK_QTY'.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
    .word_used_drw(),                             // word used quantity during write, asynchronous, minimum 0 and maximum 'BLOCK_LEN_WR * BLOCK_QTY'.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    
    .bloc_used_wr(bloc_used),                     // block used quantity, on write clock, minimum 0 and maximum BLOCK_QTY.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               
    .bloc_used_rd(bloc_used_rd),                  // block used quantity, on read clock, minimum 0 and maximum BLOCK_QTY.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                
    .bloc_used(),                                 // block used quantity, asynchronous, minimum 0 and maximum BLOCK_QTY.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 
    .bloc_full(),                                 // block full                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          
    .bloc_empty(bloc_empty),                      // block empty                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
    .overflow(),                                  // input data overflow                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 
    .underflow(),                                 // output data underflow                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               
    .data_rd_m(0),                                // memory read data                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    
    .data_wr_m({data_imag_wr_m, data_real_wr_m}), // memory write data                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
    .bloc_addr_rd_m(bloc_addr_rd_m),              // memory read block address                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           
    .base_addr_rd_m(),                            // memory read base address                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            
    .segm_addr_rd_m(),                            // memory read segment address                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
    .offs_addr_rd_m(),                            // memory read offset address                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          
    .word_addr_rd_m(word_addr_rd_m),              // memory read word address                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            
    .bloc_addr_wr_m(bloc_addr_wr_m),              // memory write block address                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          
    .base_addr_wr_m(),                            // memory write base address                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           
    .offs_addr_wr_m(),                            // memory write offset address                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
    .word_addr_wr_m(word_addr_wr_m),              // memory write word address                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           
    .en_rd_m(),                                   // memory read enable                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  
    .en_wr_m(en_wr_m),                            // memory write enable                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 
    .sop_rd_m(),                                  // memory read start of packet                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
    .sop_wr_m(sop_wr_m),                          // memory write start of packet                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        
    .eop_rd_m(eop_rd_m),                          // memory read end of packet                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           
    .eop_wr_m(eop_wr_m)                           // memory write end of packet                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          
  );                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     
           
// cpr_ram cpr_ram_real (         
//   .data(data_real_wr_m),     
//   .wraddress(word_addr_wr_m),           
//   .rdaddress(word_addr_rd_m),           
//   .wren(en_wr_m),                       
//   .wrclock(clk_wr),                     
//   .rdclock(clk_rd),                     
//   .q(dmem_real)                         
// );                                      
//                                       
// cpr_ram cpr_ram_imag (                    
//   .data(data_imag_wr_m),                
//   .wraddress(word_addr_wr_m),           
//   .rdaddress(word_addr_rd_m),           
//   .wren(en_wr_m),                       
//   .wrclock(clk_wr),                     
//   .rdclock(clk_rd),                     
//   .q(dmem_imag)                         
// );                                      
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
  cpr_ram cpr_ram_real (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
    .dina  (data_real_wr_m),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             
    .addra (word_addr_wr_m),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             
    .addrb (word_addr_rd_m),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             
    .wea   (en_wr_m),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    
    .clka  (clk_wr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     
    .clkb  (clk_rd),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     
    .doutb (dmem_real)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
  );                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
  cpr_ram cpr_ram_imag (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
    .dina (data_imag_wr_m),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
    .addra(word_addr_wr_m),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
    .addrb(word_addr_rd_m),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
    .wea  (en_wr_m),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     
    .clka (clk_wr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      
    .clkb (clk_rd),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      
    .doutb(dmem_imag)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    
  );                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
endmodule                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                